`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:48:58 11/01/2008 
// Design Name: 
// Module Name:    SP2 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module PS2(clk, rst, ps2_clk, ps2_data, data2);

input 	    clk, rst, ps2_clk , ps2_data;
output[10:0] data2;


reg [3:0] 	 i;
reg [10:0] 	 data;
reg [10:0] 	 data2;


reg [2:0] 	 ps2_clkr;
always @(posedge clk) 
	ps2_clkr <= {ps2_clkr[1:0], ps2_clk}; // ׼����ȡ�ӿڵ�ƽ�ź�

//ȷ�������غ��½���
wire ps2_clk_risingedge  = (ps2_clkr[2:1]==2'b01); 
wire ps2_clk_fallingedge = (ps2_clkr[2:1]==2'b10);


always @(posedge clk)
if(rst)
	i <= 0;
else begin
	if(ps2_clk_fallingedge)begin
		data2[i] <= data[i];   // �����һλ����
		data[i]  <= ps2_data;  //���뵱ǰ�ӿڴ�������λ
		if(i<10) 			//������ȡʮһ������λ�������굱ǰ���ݰ�
			i <= i+1;
		else 
			i <= 0;
	end
end

endmodule

